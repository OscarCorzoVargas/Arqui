module ROM #(parameter ROM_BUS_In=11, parameter ROM_BUS_Out=41)(
	//////////// OUTPUTS //////////
	ROM_DataBUS_Out,
	//////////// INPUTS //////////
	ROM_DataBUS_In
	
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
	output reg	[ROM_BUS_Out-1:0] ROM_DataBUS_Out;
	input			[ROM_BUS_In-1:0] ROM_DataBUS_In;

//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
	always@(*)
	begin
	case (ROM_DataBUS_In)	
	// Example to more outputs: WaitStart: begin sResetCounter = 0; sCuenteUP = 0; end
		11'b00000000000: ROM_DataBUS_Out = 41'b00011000001100000111010010100000000000000;//0
		11'b00000000001: ROM_DataBUS_Out = 41'b00000000000000000000000010111100000000000;//1
		
		
		//Load instructions
		11'b11100000000: ROM_DataBUS_Out = 41'b00000010000001001000000100010111100000010;//1792
		11'b11100000001: ROM_DataBUS_Out = 41'b00100000010000000000110010111011111111111;//1793
		11'b11100000010: ROM_DataBUS_Out = 41'b00011100000000001000000110000000000000000;//1794
		11'b11100000011: ROM_DataBUS_Out = 41'b00000010010000001000000100011011100000001;//1795 
//		//Storage instructions
//		11'b11100010000: ROM_DataBUS_Out = 41'b00000010000001001000000100010111100000001;//1808
//		11'b11100010001: ROM_DataBUS_Out = 41'b00011100000000000111000111111000000101000;//1809
//		11'b00000101000: ROM_DataBUS_Out = 41'b00011100000000000111000111100000000000000;//40
//		11'b00000101001: ROM_DataBUS_Out = 41'b00011100000000000111000111100000000000000;//41
//		11'b00000101010: ROM_DataBUS_Out = 41'b00011100000000100101000111100000000000000;//42
//		11'b00000101011: ROM_DataBUS_Out = 41'b10010100000000100101000111100000000000000;//43
//		11'b00000101100: ROM_DataBUS_Out = 41'b10000100000001000000001010111011111111111;//44
//		11'b11100010010: ROM_DataBUS_Out = 41'b10010100000000100001000110000000000000000;//1810
//		11'b11100010011: ROM_DataBUS_Out = 41'b00000011000010100001000100011011100010001;//1811
//		
		//ADDCC instructions
		11'b11001000000: ROM_DataBUS_Out = 41'b00000000000000000000000010110111001000010;//1600
		11'b11001000001: ROM_DataBUS_Out = 41'b00000010000001000000100001111011111111111;//1601
		11'b11001000010: ROM_DataBUS_Out = 41'b00011100000000001000000110000000000000000;//1602
		11'b11001000011: ROM_DataBUS_Out = 41'b00000010010000000000100001111011111111111;//1603
		
//		//Branch instructions
		11'b10001000000: ROM_DataBUS_Out = 41'b00000000000000000000000010111000000000010;//1088
		11'b10001011100: ROM_DataBUS_Out = 41'b00000000000000000000000010111000000000010;//1116
		11'b00000000010: ROM_DataBUS_Out = 41'b00011100000000001000000101000000000000000;//2
		11'b00000000011: ROM_DataBUS_Out = 41'b00100000000000001000000111100000000000000;//3 
		11'b00000000100: ROM_DataBUS_Out = 41'b00100000000000001000000111100000000000000;//4 
		11'b00000000101: ROM_DataBUS_Out = 41'b00011100000000000111000111100000000000000;//5 
		11'b00000000110: ROM_DataBUS_Out = 41'b00011100000000000111000111100000000000000;//6 
		11'b00000000111: ROM_DataBUS_Out = 41'b00011100000000000111000111100000000000000;//7 
		11'b00000001000: ROM_DataBUS_Out = 41'b00011100001110000111000100010100000001100;// preguntar //8
		11'b00000001001: ROM_DataBUS_Out = 41'b00011100001110000111000100010100000001101;// preguntar //9
		11'b00000001010: ROM_DataBUS_Out = 41'b00011100001110000111000100001000000001100;// preguntar //10
		11'b00000001011: ROM_DataBUS_Out = 41'b00000000000000000000000010111011111111111;//11 
		11'b00000001100: ROM_DataBUS_Out = 41'b00011000010000000110000100011000000000000;//12 
		11'b00000001101: ROM_DataBUS_Out = 41'b00011100001110000111000100010100000010000;//13 
		11'b00000001110: ROM_DataBUS_Out = 41'b00000000000000000000000010110000000001100;//14 
		11'b00000001111: ROM_DataBUS_Out = 41'b00000000000000000000000010111011111111111;//15 
		11'b00000010000: ROM_DataBUS_Out = 41'b00000000000000000000000010110100000010011;//16 
		11'b00000010001: ROM_DataBUS_Out = 41'b00000000000000000000000010100100000001100;//17 
		11'b00000010010: ROM_DataBUS_Out = 41'b00000000000000000000000010111011111111111;//18 
		11'b00000010011: ROM_DataBUS_Out = 41'b00000000000000000000000010101100000001100;//19 
		11'b00000010100: ROM_DataBUS_Out = 41'b00000000000000000000000010111011111111111;//20 
		11'b11111111111: ROM_DataBUS_Out = 41'b00011000000000000110000111011000000000000;//2047

		
//		//


		default :   ROM_DataBUS_Out = 41'b00011000001100000111010010100000000000000; // channel 0 is selected 
		endcase
	end
//=======================================================
//  Outputs
//=======================================================
// OUTPUT LOGIC : COMBINATIONAL

endmodule
